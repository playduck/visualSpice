.title Gleichrichter
.model filesrc filesource (file="__INPUT_FILE__" amploffset=[0] amplscale=[0.0005]
+                           timeoffset=0 timescale=1
+                           timerelative=false amplstep=false)

.model ads1 sidiode(Roff=1000 Ron=0.7 Rrev=0.2 Vfwd=1
+       Vrev=10 Revepsilon=0.2 Epsilon=0.2 Ilimit=7 Revilimit=15)

a1 %vd([input, b]) filesrc

ad1 input out ads1
ad2 0 input ads1
ad3 0 b ads1
ad4 b out ads1

R1 out 0 10k
C1 out 0 100e-6

.tran 100u 5
.save all
.end
