.title Basic low pass filter circuit

.control
** uncomment to save as ascii file
* set wr_singlescale
* set wr_vecnames
* tran 80u 4
* wrdata __OUTPUT_FILE__ V(input) V(2)
.endc

.model filesrc filesource (file="__INPUT_FILE__" amploffset=[0] amplscale=[1]
+                           timeoffset=0 timescale=1
+                           timerelative=false amplstep=false)

a1 %v([input]) filesrc

R1 input 1 1k
L1 1 2 2.2m
C1 2 0 24e-6
R2 2 0 1k

.tran 80u 4
.save all
.end
